library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity Multiplexer_2_to_1 is
port (	-- Datenleitungen
		A: in STD_LOGIC; -- Eingang 1
		B: in STD_LOGIC; -- Eingang 2
		Y: out STD_LOGIC; --Ausgang
		-- Steuerleitungen
		S: in STD_LOGIC);
end Multiplexer_2_to_1;

architecture Behavior of Multiplexer_2_to_1 is
begin
	Y <= 	A when (S = '0') else
			B when (S = '1');
end Behavior;

	-- 2-zu-1 Multiplexer
	component Multiplexer_2_to_1
		port (	A, B: in STD_LOGIC;
				Y: out STD_LOGIC;
				S: in STD_LOGIC);
	end component Multiplexer_2_to_1;